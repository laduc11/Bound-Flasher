module bound_flasher (flick, clk, rst, led);
  input wire flick;
  input wire clk;
  input wire rst;
  output reg [15:0] led;
  
  reg [2:0] state;
  reg [2:0] real_state;
  reg [15:0] temp_led;
  
  reg flickFlag;
  
  //FLIP FLOP OUTPUT
  always @(posedge clk or negedge rst) begin
    if (rst == 1'b0) begin
      led <= 16'b0;
    end
    else begin
      led <= temp_led;
    end
  end
  
  always @(state or led) begin
    if (state == 3'b0) begin
      temp_led = 16'b0;
    end
    else if (state == 3'b001 || state == 3'b011 || state == 3'b101) begin
      temp_led = (led << 1) | 1;
    end
    else if (state == 3'b010 || state == 3'b100 || state == 3'b110) begin
      temp_led = led >> 1;
    end
    else begin
      temp_led = 16'b0;
    end
  end
  
  //FLIP FLOP STATE
  always @(posedge clk or negedge rst) begin
    if (rst == 1'b0) begin
      real_state <= 3'b0;
    end
    else begin
      real_state <= state;
    end
  end
  
  always @(flick or real_state or led or rst) begin
    if (rst == 1'b0) begin
      state = 3'b0;
    end
    else begin
    case (real_state)
      3'b0: begin
        if (flick == 1) begin
          state = 3'b001;
        end
      end
      
      3'b001: begin
        if (led[15] == 1) begin
          state = 3'b010;
        end
      end
      
      3'b010: begin	// state 2
        if (flick == 1 && led[5] == 0) begin
          state = 3'b001;
        end
        else if (led[5] == 0 && flickFlag == 0) begin
          state = 3'b011;
        end
      end
      
      3'b011: begin
        if (led[10] == 1) begin
          state = 3'b100;
        end
      end
      
      3'b100: begin	// state 4
        if (flick == 1 && led[5:4] == 2'b01) begin
          state = 3'b011;
        end
        else if (flick == 1 && led[0] == 0) begin
          state = 3'b011;
        end  
        else if (led[0] == 0 && flickFlag == 0) begin
          state = 3'b101;
        end
      end
      
      3'b101: begin
        if (led[5] == 1) begin
          state = 3'b110;
        end
      end
      
      3'b110: begin
        if (led[0] == 0) begin
          state = 3'b000;
        end
      end
      
      default: state = 3'b000;
    endcase
    end
  end
  
  always @(flick or rst or real_state or led) begin
    if (rst == 1'b0) begin
      flickFlag = 1'b0;
    end
    else if (flick == 1'b1 && real_state == 3'b010 && led[5] == 0) begin
      flickFlag = 1'b1;
    end
    else if (flick == 1'b1 && real_state == 3'b100 && led[5:4] == 2'b01) begin
      flickFlag = 1'b1;
    end    
    else if (flick == 1'b1 && real_state == 3'b100 && led[0] == 0) begin
      flickFlag = 1'b1;
    end 
    else if (led[5] == 1) begin
      flickFlag = 1'b0;
    end
    else if (real_state == 3'b011 && led[1:0] == 2'b01) begin
      flickFlag = 1'b0;
    end
  end

endmodule
